module COMP64 (x_a, x_b, wx);
  input  [63:0] x_a, x_b;
  output wx;
  wire [63:0] XOR;
  wire [31:0] temp;
  wire GT2_32,GT2_31,GT2_30,GT2_29,GT2_28,GT2_27,GT2_26,GT2_25,GT2_24,GT2_23,GT2_22,GT2_21,GT2_20,GT2_19,GT2_18,GT2_17;
  wire GT2_16,GT2_15,GT2_14,GT2_13,GT2_12,GT2_11,GT2_10,GT2_9,GT2_8,GT2_7,GT2_6,GT2_5,GT2_4,GT2_3,GT2_2,GT2_1;
  wire GT4_16,GT4_15,GT4_14,GT4_13,GT4_12,GT4_11,GT4_10,GT4_9,GT4_8,GT4_7,GT4_6,GT4_5,GT4_4,GT4_3,GT4_2,GT4_1;
  wire GT8_8,GT8_7,GT8_6,GT8_5,GT8_4,GT8_3,GT8_2,GT8_1;
  wire GT16_4,GT16_3,GT16_2,GT16_1;
  wire GT32_1,GT32_2;
  wire GT64_1;
  wire AND63_60,AND55_52,AND47_44,AND39_36,AND31_28,AND23_20,AND15_12,AND59_56,AND63_56,AND43_40,AND51_48,AND35_32,AND63_32,AND19_16,AND27_24,AND31_16,AND11_8,AND7_4,AND31_24; 
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[63]= x_a[63] ^ (!x_b[63]);
  assign XOR[62]= x_a[62] ^ (!x_b[62]);
  assign GT2_32 = (x_a[63] & (!x_b[63])) ^ (XOR[63] & x_a[62] & (!x_b[62]));//depth1
 
  assign XOR[61] = x_a[61] ^ (!x_b[61]);
  assign XOR[60] = x_a[60] ^ (!x_b[60]);
  assign GT2_31 = (x_a[61] & (!x_b[61])) ^ (XOR[61] & x_a[60] & (!x_b[60]));//depth1
  
  assign temp[16] = XOR[63] & XOR[62] & GT2_31;//depth2
  assign GT4_16 = temp[16] ^ GT2_32;//depth2 
  /////////////////////////////////////////////
  assign XOR[59]= x_a[59] ^ (!x_b[59]);
  assign XOR[58]= x_a[58] ^ (!x_b[58]);
  assign GT2_30 = (x_a[59] & (!x_b[59])) ^ (XOR[59] & x_a[58] & (!x_b[58]));//depth1
 
  assign XOR[57] = x_a[57] ^ (!x_b[57]);
  assign XOR[56] = x_a[56] ^ (!x_b[56]);
  assign GT2_29 = (x_a[57] & (!x_b[57])) ^ (XOR[57] & x_a[56] & (!x_b[56]));//depth1
  
  //assign temp[15] = XOR[59] & XOR[58] & GT2_29;//depth2
  //assign GT4_15 = temp[15] ^ GT2_30;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[24]= XOR[63] & XOR[62] & XOR[61] & XOR[60];//depth1
  assign AND63_60= (temp[24] & GT2_30) ^ (temp[24] & XOR[59] & XOR[58] & GT2_29);//depth2
  assign GT8_8 = AND63_60 ^ GT4_16;
   /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[55]= x_a[55] ^ (!x_b[55]);
  assign XOR[54]= x_a[54] ^ (!x_b[54]);
  assign GT2_28 = (x_a[55] & (!x_b[55])) ^ (XOR[55] & x_a[54] & (!x_b[54]));//depth1
 
  assign XOR[53] = x_a[53] ^ (!x_b[53]);
  assign XOR[52] = x_a[52] ^ (!x_b[52]);
  assign GT2_27 = (x_a[53] & (!x_b[53])) ^ (XOR[53] & x_a[52] & (!x_b[52]));//depth1
  
  assign temp[14] = XOR[55] & XOR[54] & GT2_27;//depth2
  assign GT4_14 = temp[14] ^ GT2_28;//depth2 
  /////////////////////////////////////////////
  assign XOR[51]= x_a[51] ^ (!x_b[51]);
  assign XOR[50]= x_a[50] ^ (!x_b[50]);
  assign GT2_26 = (x_a[51] & (!x_b[51])) ^ (XOR[51] & x_a[50] & (!x_b[50]));//depth1
 
  assign XOR[49] = x_a[49] ^ (!x_b[49]);
  assign XOR[48] = x_a[48] ^ (!x_b[48]);
  assign GT2_25 = (x_a[49] & (!x_b[49])) ^ (XOR[49] & x_a[48] & (!x_b[48]));//depth1
  
  //assign temp[13] = XOR[51] & XOR[50] & GT2_25;//depth2
  //assign GT4_13 = temp[13] ^ GT2_26;//depth2
   /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[23]= XOR[55] & XOR[54] & XOR[53] & XOR[52];//depth1
  assign AND55_52= (temp[23] & GT2_26) ^ (temp[23] & XOR[51] & XOR[50] & GT2_25);//depth2
  assign GT8_7 = AND55_52 ^ GT4_14;
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign AND59_56= XOR[59] & XOR[58] & XOR[57] & XOR[56];//depth1
  assign temp[28]= AND59_56& temp[24];//depth2
  assign AND63_56=temp[28]&GT8_7;//depth3
  assign GT16_4 = AND63_56 ^ GT8_8;//depth3
  /////////////////////////////////////////////
  /////////////////////////////////////////////
  ////////////////////////////////////////////
  
  assign XOR[47]= x_a[47] ^ (!x_b[47]);
  assign XOR[46]= x_a[46] ^ (!x_b[46]);
  assign GT2_24 = (x_a[47] & (!x_b[47])) ^ (XOR[47] & x_a[46] & (!x_b[46]));//depth1
 
  assign XOR[45] = x_a[45] ^ (!x_b[45]);
  assign XOR[44] = x_a[44] ^ (!x_b[44]);
  assign GT2_23 = (x_a[45] & (!x_b[45])) ^ (XOR[45] & x_a[44] & (!x_b[44]));//depth1
  
  assign temp[12] = XOR[47] & XOR[46] & GT2_23;//depth2
  assign GT4_12 = temp[12] ^ GT2_24;//depth2
  /////////////////////////////////////////////
  assign XOR[43]= x_a[43] ^ (!x_b[43]);
  assign XOR[42]= x_a[42] ^ (!x_b[42]);
  assign GT2_22 = (x_a[43] & (!x_b[43])) ^ (XOR[43] & x_a[42] & (!x_b[42]));//depth1
 
  assign XOR[41] = x_a[41] ^ (!x_b[41]);
  assign XOR[40] = x_a[40] ^ (!x_b[40]);
  assign GT2_21 = (x_a[41] & (!x_b[41])) ^ (XOR[41] & x_a[40] & (!x_b[40]));//depth1
  
  //assign temp[11] = XOR[43] & XOR[42] & GT2_21;//depth2
  //assign GT4_11 = temp[11] ^ GT2_22;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[22]= XOR[47] & XOR[46] & XOR[45] & XOR[44];//depth1
  assign AND47_44= (temp[22] & GT2_22) ^ (temp[22] & XOR[43] & XOR[42] & GT2_21);//depth2
  assign GT8_6 = AND47_44 ^ GT4_12;
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[39]= x_a[39] ^ (!x_b[39]);
  assign XOR[38]= x_a[38] ^ (!x_b[38]);
  assign GT2_20 = (x_a[39] & (!x_b[39])) ^ (XOR[39] & x_a[38] & (!x_b[38]));//depth1
 
  assign XOR[37] = x_a[37] ^ (!x_b[37]);
  assign XOR[36] = x_a[36] ^ (!x_b[36]);
  assign GT2_19 = (x_a[37] & (!x_b[37])) ^ (XOR[37] & x_a[36] & (!x_b[36]));//depth1
  
  assign temp[10] = XOR[39] & XOR[38] & GT2_19;//depth2
  assign GT4_10 = temp[10] ^ GT2_20;//depth2
  ///////////////////////////////////////////// 
  assign XOR[35]= x_a[35] ^ (!x_b[35]);
  assign XOR[34]= x_a[34] ^ (!x_b[34]);
  assign GT2_18 = (x_a[35] & (!x_b[35])) ^ (XOR[35] & x_a[34] & (!x_b[34]));//depth1
 
  assign XOR[33] = x_a[33] ^ (!x_b[33]);
  assign XOR[32] = x_a[32] ^ (!x_b[32]);
  assign GT2_17 = (x_a[33] & (!x_b[33])) ^ (XOR[33] & x_a[32] & (!x_b[32]));//depth1
  
  //assign temp[9] = XOR[35] & XOR[34] & GT2_17;//depth2
 // assign GT4_9 = temp[9] ^ GT2_18;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[21]= XOR[39] & XOR[38] & XOR[37] & XOR[36];//depth1
  assign AND39_36= (temp[21] & GT2_18) ^ (temp[21] & XOR[35] & XOR[34] & GT2_17);//depth2
  assign GT8_5 = AND39_36 ^ GT4_10;
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign AND43_40= XOR[43] & XOR[42] & XOR[41] & XOR[40];//depth1
  assign temp[27]= AND43_40& temp[22];//depth2
  //assign XOR47_40=temp[27]&GT8_5;//depth3
  //assign GT16_3 = XOR47_40 ^ GT8_6;//depth3
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign AND51_48= XOR[51] & XOR[50] & XOR[49] & XOR[48];//depth1
  assign temp[30]= AND51_48& AND59_56& temp[24]&temp[23];//depth2
  assign AND63_32= (temp[30]&temp[27]&GT8_5) ^ (temp[30]& GT8_6);//depth3
  assign GT32_2 = AND63_32 ^ GT16_4;//depth3
  /////////////////////////////////////////////
  /////////////////////////////////////////////
  /////////////////////////////////////////////
  assign XOR[31]= x_a[31] ^ (!x_b[31]);
  assign XOR[30]= x_a[30] ^ (!x_b[30]);
  assign GT2_16 = (x_a[31] & (!x_b[31])) ^ (XOR[31] & x_a[30] & (!x_b[30]));//depth1
 
  assign XOR[29] = x_a[29] ^ (!x_b[29]);
  assign XOR[28] = x_a[28] ^ (!x_b[28]);
  assign GT2_15 = (x_a[29] & (!x_b[29])) ^ (XOR[29] & x_a[28] & (!x_b[28]));//depth1
  
  assign temp[8] = XOR[31] & XOR[30] & GT2_15;//depth2
  assign GT4_8 = temp[8] ^ GT2_16;//depth2
  ///////////////////////////////////////////// 
  assign XOR[27]= x_a[27] ^ (!x_b[27]);
  assign XOR[26]= x_a[26] ^ (!x_b[26]);
  assign GT2_14 = (x_a[27] & (!x_b[27])) ^ (XOR[27] & x_a[26] & (!x_b[26]));//depth1
 
  assign XOR[25] = x_a[25] ^ (!x_b[25]);
  assign XOR[24] = x_a[24] ^ (!x_b[24]);
  assign GT2_13 = (x_a[25] & (!x_b[25])) ^ (XOR[25] & x_a[24] & (!x_b[24]));//depth1
  
  //assign temp[7] = XOR[27] & XOR[26] & GT2_13;//depth2
  //assign GT4_7 = temp[7] ^ GT2_14;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[20]= XOR[31] & XOR[30] & XOR[29] & XOR[28];//depth1
  assign AND31_28= (temp[20] & GT2_14) ^ (temp[20] & XOR[27] & XOR[26] & GT2_13);//depth2
  assign GT8_4 = AND31_28 ^ GT4_8;
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[23]= x_a[23] ^ (!x_b[23]);
  assign XOR[22]= x_a[22] ^ (!x_b[22]);
  assign GT2_12 = (x_a[23] & (!x_b[23])) ^ (XOR[23] & x_a[22] & (!x_b[22])); //depth1
 
  assign XOR[21] = x_a[21] ^ (!x_b[21]);
  assign XOR[20] = x_a[20] ^ (!x_b[20]);
  assign GT2_11 = (x_a[21] & (!x_b[21])) ^ (XOR[21] & x_a[20] & (!x_b[20])); //depth1
  
  assign temp[6] = XOR[23] & XOR[22] & GT2_11;//depth2
  assign GT4_6 = temp[6] ^ GT2_12;//depth2
  ///////////////////////////////////////////// 
  assign XOR[19]= x_a[19] ^ (!x_b[19]);
  assign XOR[18]= x_a[18] ^ (!x_b[18]);
  assign GT2_10 = (x_a[19] & (!x_b[19])) ^ (XOR[19] & x_a[18] & (!x_b[18]));//depth1
 
  assign XOR[17] = x_a[17] ^ (!x_b[17]);
  assign XOR[16] = x_a[16] ^ (!x_b[16]);
  assign GT2_9 = (x_a[17] & (!x_b[17])) ^ (XOR[17] & x_a[16] & (!x_b[16]));//depth1
  
  //assign temp[5] = XOR[19] & XOR[18] & GT2_9;//depth2
  //assign GT4_5 = temp[5] ^ GT2_10;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[19]= XOR[23] & XOR[22] & XOR[21] & XOR[20];//depth1
  assign AND23_20= (temp[19] & GT2_10) ^ (temp[19] & XOR[19] & XOR[18] & GT2_9);//depth2
  assign GT8_3 = AND23_20 ^ GT4_6;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign AND27_24= XOR[27] & XOR[26] & XOR[25] & XOR[24];//depth1
  assign temp[26]= AND27_24& temp[20];//depth2
  assign AND31_24=temp[26]&GT8_3;//depth3
  assign GT16_2 = AND31_24 ^ GT8_4;//depth3
  /////////////////////////////////////////////
  /////////////////////////////////////////////
  ////////////////////////////////////////////
  assign XOR[15]= x_a[15] ^ (!x_b[15]); //depth1
  assign XOR[14]= x_a[14] ^ (!x_b[14]);
  assign GT2_8 = (x_a[15] & (!x_b[15])) ^ (XOR[15] & x_a[14] & (!x_b[14]));//depth1
 
  assign XOR[13] = x_a[13] ^ (!x_b[13]);
  assign XOR[12] = x_a[12] ^ (!x_b[12]);
  assign GT2_7 = (x_a[13] & (!x_b[13])) ^ (XOR[13] & x_a[12] & (!x_b[12]));//depth1
  
  assign temp[4] = XOR[15] & XOR[14] & GT2_7;//depth2
  assign GT4_4 = temp[4] ^ GT2_8;//depth2
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[11]= x_a[11] ^ (!x_b[11]);
  assign XOR[10]= x_a[10] ^ (!x_b[10]);
  assign GT2_6 = (x_a[11] & (!x_b[11])) ^ (XOR[11] & x_a[10] & (!x_b[10]));//depth1
 
  assign XOR[9] = x_a[9] ^ (!x_b[9]);
  assign XOR[8] = x_a[8] ^ (!x_b[8]);
  assign GT2_5 = (x_a[9] & (!x_b[9])) ^ (XOR[9] & x_a[8] & (!x_b[8]));//depth1
  
  //assign temp[3] = XOR[11] & XOR[10] & GT2_5;//depth2
  //assign GT4_3 = temp[3] ^ GT2_6;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[18]= XOR[15] & XOR[14] & XOR[13] & XOR[12];//depth1
  assign AND15_12= (temp[18] & GT2_6) ^ (temp[18] & XOR[11] & XOR[10] & GT2_5);//depth2
  assign GT8_2 = AND15_12 ^ GT4_4;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[7]= x_a[7] ^ (!x_b[7]);
  assign XOR[6]= x_a[6] ^ (!x_b[6]);
  assign GT2_4 = (x_a[7] & (!x_b[7])) ^ (XOR[7] & x_a[6] & (!x_b[6]));//depth1
 
  assign XOR[5] = x_a[5] ^ (!x_b[5]);
  assign XOR[4] = x_a[4] ^ (!x_b[4]);
  assign GT2_3  = (x_a[5] & (!x_b[5])) ^ (XOR[5] & x_a[4] & (!x_b[4]));//depth1
  
  assign temp[2] = XOR[7] & XOR[6] & GT2_3;//depth2
  assign GT4_2 = temp[2] ^ GT2_4;//depth2
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[3]= x_a[3] ^ (!x_b[3]);
  assign XOR[2]= x_a[2] ^ (!x_b[2]);
  assign GT2_2 = (x_a[3] & (!x_b[3])) ^ (XOR[3] & x_a[2] & (!x_b[2]));//depth1
 
  assign XOR[1] = x_a[1] ^ (!x_b[1]);
  assign XOR[0] = x_a[0] ^ (!x_b[0]);
  assign GT2_1  = (x_a[1] & (!x_b[1])) ^ (XOR[1] & x_a[0] & (!x_b[0]));//depth1
  
  //assign temp[1] = XOR[3] & XOR[2] & GT2_1;//depth2
  //assign GT4_1 = temp[1] ^ GT2_2;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[17]= XOR[7] & XOR[6] & XOR[5] & XOR[4];//depth1
  assign AND7_4= (temp[17] & GT2_2) ^ (temp[17] & XOR[3] & XOR[2] & GT2_1);//depth2
  assign GT8_1 = AND7_4 ^ GT4_2;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign AND11_8= XOR[11] & XOR[10] & XOR[9] & XOR[8];//depth1
  assign temp[25]= AND11_8& temp[18];//depth2
  //assign XOR15_8=temp[25]&GT8_1;//depth3
  //assign GT16_1 = XOR15_8 ^ GT8_2;//depth3
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign AND19_16= XOR[19] & XOR[18] & XOR[17] & XOR[16];//depth1
  assign temp[29]= AND19_16& AND27_24& temp[20]&temp[19];//depth2
  assign AND31_16= (temp[29]&temp[25]&GT8_1) ^ (temp[29]& GT8_2);//depth3
  assign GT32_1 = AND31_16 ^ GT16_2;//depth3
   /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign AND35_32= XOR[35] & XOR[34] & XOR[33] & XOR[32];//depth1
  assign temp[31]= (temp[24] & temp[23] & temp[22] & temp[21]) & (AND35_32& AND43_40& AND51_48& AND59_56);//depth2
  assign AND63_32= (temp[31]&GT32_1);//depth4
  assign GT64_1 = AND63_32 ^ GT32_2;//depth4
  /////////////////////////////////////////////
  /////////////////////////////////////////////
  ///////////////////////////////////////////// 
  assign wx = GT64_1;
endmodule



