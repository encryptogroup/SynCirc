module __f32sub__main(
  input wire [31:0] x,
  input wire [31:0] y,
  output wire [31:0] out
);
  wire [7:0] y_bexp__4;
  wire [7:0] x_bexp__4;
  wire [8:0] sum;
  wire [22:0] tuple_index_1846;
  wire [22:0] y_fraction__4;
  wire [7:0] y_bexp__5;
  wire [22:0] y_fraction__5;
  wire [7:0] incremented_sum__1;
  wire [27:0] wide_y;
  wire [7:0] x_bexpbs_difference__2;
  wire [7:0] x_bexp__5;
  wire [27:0] wide_y__1;
  wire [7:0] sub_1865;
  wire [22:0] x_fraction__1;
  wire [27:0] dropped;
  wire y_sign__2;
  wire [27:0] wide_x;
  wire tuple_index_1877;
  wire [27:0] wide_x__1;
  wire x_sign__1;
  wire y_sign__3;
  wire [27:0] neg_1883;
  wire [27:0] sticky;
  wire [27:0] xddend_y__1;
  wire [24:0] sel_1890;
  wire [25:0] add_1895;
  wire [27:0] concat_1898;
  wire [27:0] xbs_fraction__1;
  wire [27:0] reverse_1902;
  wire [28:0] one_hot_1903;
  wire [4:0] encode_1904;
  wire cancel__2;
  wire carry_bit;
  wire [27:0] leading_zeroes;
  wire [26:0] carry_fraction;
  wire [27:0] add_1921;
  wire [2:0] concat_1922;
  wire [26:0] carry_fraction__1;
  wire [26:0] cancel_fraction;
  wire [26:0] shifted_fraction;
  wire [2:0] normal_chunk;
  wire [2:0] fraction_shift__3;
  wire [1:0] half_way_chunk;
  wire [24:0] add_1937;
  wire do_round_up;
  wire [27:0] rounded_fraction;
  wire rounding_carry;
  wire [8:0] add_1948;
  wire [9:0] add_1956;
  wire [9:0] wide_exponent;
  wire [9:0] wide_exponent__1;
  wire [7:0] MAX_EXPONENT;
  wire [7:0] MAX_EXPONENT__1;
  wire [8:0] wide_exponent__2;
  wire [7:0] MAX_EXPONENT__3;
  wire [7:0] MAX_EXPONENT__4;
  wire eq_1977;
  wire eq_1978;
  wire eq_1979;
  wire eq_1980;
  wire ne_1983;
  wire ne_1985;
  wire fraction_is_zero;
  wire [2:0] fraction_shift__2;
  wire [2:0] fraction_shift__4;
  wire is_operand_inf;
  wire and_reduce_2002;
  wire has_pos_inf;
  wire has_neg_inf;
  wire [2:0] fraction_shift__1;
  wire [2:0] concat_2012;
  wire [27:0] shrl_2015;
  wire is_result_nan;
  wire result_sign;
  wire [22:0] result_fraction;
  wire result_sign__1;
  wire [7:0] MAX_EXPONENT__2;
  wire [22:0] result_fraction__3;
  wire [22:0] FRACTION_HIGH_BIT;
  wire result_sign__2;
  wire [7:0] result_exponent__2;
  wire [22:0] result_fraction__4;
  assign y_bexp__4 = y[30:23];
  assign x_bexp__4 = x[30:23];
  assign sum = {1'h0, x_bexp__4} + {1'h0, ~y_bexp__4};
  assign tuple_index_1846 = x[22:0];
  assign y_fraction__4 = y[22:0];
  assign y_bexp__5 = sum[8] ? y_bexp__4 : x_bexp__4;
  assign y_fraction__5 = sum[8] ? y_fraction__4 : tuple_index_1846;
  assign incremented_sum__1 = sum[7:0] + 8'h01;
  assign wide_y = {2'h1, y_fraction__5, 3'h0};
  assign x_bexpbs_difference__2 = sum[8] ? incremented_sum__1 : ~sum[7:0];
  assign x_bexp__5 = sum[8] ? x_bexp__4 : y_bexp__4;
  assign wide_y__1 = wide_y & {28{y_bexp__5 != 8'h00}};
  assign sub_1865 = 8'h1c - x_bexpbs_difference__2;
  assign x_fraction__1 = sum[8] ? tuple_index_1846 : y_fraction__4;
  assign dropped = sub_1865 >= 8'h1c ? 28'h000_0000 : wide_y__1 << sub_1865;
  assign y_sign__2 = y[31:31];
  assign wide_x = {2'h1, x_fraction__1, 3'h0};
  assign tuple_index_1877 = x[31:31];
  assign wide_x__1 = wide_x & {28{x_bexp__5 != 8'h00}};
  assign x_sign__1 = sum[8] ? tuple_index_1877 : ~y_sign__2;
  assign y_sign__3 = sum[8] ? ~y_sign__2 : tuple_index_1877;
  assign neg_1883 = -wide_x__1;
  assign sticky = {27'h000_0000, dropped[27:3] != 25'h000_0000};
  assign xddend_y__1 = (x_bexpbs_difference__2 >= 8'h1c ? 28'h000_0000 : wide_y__1 >> x_bexpbs_difference__2) | sticky;
  assign sel_1890 = x_sign__1 ^ y_sign__3 ? neg_1883[27:3] : wide_x__1[27:3];
  assign add_1895 = {{1{sel_1890[24]}}, sel_1890} + {1'h0, xddend_y__1[27:3]};
  assign concat_1898 = {add_1895[24:0], xddend_y__1[2:0]};
  assign xbs_fraction__1 = add_1895[25] ? -concat_1898 : concat_1898;
  assign reverse_1902 = {xbs_fraction__1[0], xbs_fraction__1[1], xbs_fraction__1[2], xbs_fraction__1[3], xbs_fraction__1[4], xbs_fraction__1[5], xbs_fraction__1[6], xbs_fraction__1[7], xbs_fraction__1[8], xbs_fraction__1[9], xbs_fraction__1[10], xbs_fraction__1[11], xbs_fraction__1[12], xbs_fraction__1[13], xbs_fraction__1[14], xbs_fraction__1[15], xbs_fraction__1[16], xbs_fraction__1[17], xbs_fraction__1[18], xbs_fraction__1[19], xbs_fraction__1[20], xbs_fraction__1[21], xbs_fraction__1[22], xbs_fraction__1[23], xbs_fraction__1[24], xbs_fraction__1[25], xbs_fraction__1[26], xbs_fraction__1[27]};
  assign one_hot_1903 = {reverse_1902[27:0] == 28'h000_0000, reverse_1902[27] && reverse_1902[26:0] == 27'h000_0000, reverse_1902[26] && reverse_1902[25:0] == 26'h000_0000, reverse_1902[25] && reverse_1902[24:0] == 25'h000_0000, reverse_1902[24] && reverse_1902[23:0] == 24'h00_0000, reverse_1902[23] && reverse_1902[22:0] == 23'h00_0000, reverse_1902[22] && reverse_1902[21:0] == 22'h00_0000, reverse_1902[21] && reverse_1902[20:0] == 21'h00_0000, reverse_1902[20] && reverse_1902[19:0] == 20'h0_0000, reverse_1902[19] && reverse_1902[18:0] == 19'h0_0000, reverse_1902[18] && reverse_1902[17:0] == 18'h0_0000, reverse_1902[17] && reverse_1902[16:0] == 17'h0_0000, reverse_1902[16] && reverse_1902[15:0] == 16'h0000, reverse_1902[15] && reverse_1902[14:0] == 15'h0000, reverse_1902[14] && reverse_1902[13:0] == 14'h0000, reverse_1902[13] && reverse_1902[12:0] == 13'h0000, reverse_1902[12] && reverse_1902[11:0] == 12'h000, reverse_1902[11] && reverse_1902[10:0] == 11'h000, reverse_1902[10] && reverse_1902[9:0] == 10'h000, reverse_1902[9] && reverse_1902[8:0] == 9'h000, reverse_1902[8] && reverse_1902[7:0] == 8'h00, reverse_1902[7] && reverse_1902[6:0] == 7'h00, reverse_1902[6] && reverse_1902[5:0] == 6'h00, reverse_1902[5] && reverse_1902[4:0] == 5'h00, reverse_1902[4] && reverse_1902[3:0] == 4'h0, reverse_1902[3] && reverse_1902[2:0] == 3'h0, reverse_1902[2] && reverse_1902[1:0] == 2'h0, reverse_1902[1] && !reverse_1902[0], reverse_1902[0]};
  assign encode_1904 = {one_hot_1903[16] | one_hot_1903[17] | one_hot_1903[18] | one_hot_1903[19] | one_hot_1903[20] | one_hot_1903[21] | one_hot_1903[22] | one_hot_1903[23] | one_hot_1903[24] | one_hot_1903[25] | one_hot_1903[26] | one_hot_1903[27] | one_hot_1903[28], one_hot_1903[8] | one_hot_1903[9] | one_hot_1903[10] | one_hot_1903[11] | one_hot_1903[12] | one_hot_1903[13] | one_hot_1903[14] | one_hot_1903[15] | one_hot_1903[24] | one_hot_1903[25] | one_hot_1903[26] | one_hot_1903[27] | one_hot_1903[28], one_hot_1903[4] | one_hot_1903[5] | one_hot_1903[6] | one_hot_1903[7] | one_hot_1903[12] | one_hot_1903[13] | one_hot_1903[14] | one_hot_1903[15] | one_hot_1903[20] | one_hot_1903[21] | one_hot_1903[22] | one_hot_1903[23] | one_hot_1903[28], one_hot_1903[2] | one_hot_1903[3] | one_hot_1903[6] | one_hot_1903[7] | one_hot_1903[10] | one_hot_1903[11] | one_hot_1903[14] | one_hot_1903[15] | one_hot_1903[18] | one_hot_1903[19] | one_hot_1903[22] | one_hot_1903[23] | one_hot_1903[26] | one_hot_1903[27], one_hot_1903[1] | one_hot_1903[3] | one_hot_1903[5] | one_hot_1903[7] | one_hot_1903[9] | one_hot_1903[11] | one_hot_1903[13] | one_hot_1903[15] | one_hot_1903[17] | one_hot_1903[19] | one_hot_1903[21] | one_hot_1903[23] | one_hot_1903[25] | one_hot_1903[27]};
  assign cancel__2 = |encode_1904[4:1];
  assign carry_bit = xbs_fraction__1[27];
  assign leading_zeroes = {23'h00_0000, encode_1904};
  assign carry_fraction = xbs_fraction__1[27:1];
  assign add_1921 = leading_zeroes + 28'hfff_ffff;
  assign concat_1922 = {~(carry_bit | cancel__2), ~(carry_bit | ~cancel__2), ~(~carry_bit | cancel__2)};
  assign carry_fraction__1 = carry_fraction | {26'h000_0000, xbs_fraction__1[0]};
  assign cancel_fraction = add_1921 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__1[26:0] << add_1921;
  assign shifted_fraction = carry_fraction__1 & {27{concat_1922[0]}} | cancel_fraction & {27{concat_1922[1]}} | xbs_fraction__1[26:0] & {27{concat_1922[2]}};
  assign normal_chunk = shifted_fraction[2:0];
  assign fraction_shift__3 = 3'h4;
  assign half_way_chunk = shifted_fraction[3:2];
  assign add_1937 = {1'h0, shifted_fraction[26:3]} + 25'h000_0001;
  assign do_round_up = normal_chunk > fraction_shift__3 | half_way_chunk == 2'h3;
  assign rounded_fraction = do_round_up ? {add_1937, normal_chunk} : {1'h0, shifted_fraction};
  assign rounding_carry = rounded_fraction[27];
  assign add_1948 = {1'h0, x_bexp__5} + {8'h00, rounding_carry};
  assign add_1956 = {1'h0, add_1948} + 10'h001;
  assign wide_exponent = add_1956 - {5'h00, encode_1904};
  assign wide_exponent__1 = wide_exponent & {10{add_1895 != 26'h000_0000 | xddend_y__1[2:0] != 3'h0}};
  assign MAX_EXPONENT = 8'hff;
  assign MAX_EXPONENT__1 = 8'hff;
  assign wide_exponent__2 = wide_exponent__1[8:0] & {9{~wide_exponent__1[9]}};
  assign MAX_EXPONENT__3 = 8'hff;
  assign MAX_EXPONENT__4 = 8'hff;
  assign eq_1977 = x_bexp__5 == MAX_EXPONENT;
  assign eq_1978 = x_fraction__1 == 23'h00_0000;
  assign eq_1979 = y_bexp__5 == MAX_EXPONENT__1;
  assign eq_1980 = y_fraction__5 == 23'h00_0000;
  assign ne_1983 = x_fraction__1 != 23'h00_0000;
  assign ne_1985 = y_fraction__5 != 23'h00_0000;
  assign fraction_is_zero = add_1895 == 26'h000_0000 & xddend_y__1[2:0] == 3'h0;
  assign fraction_shift__2 = 3'h3;
  assign fraction_shift__4 = 3'h4;
  assign is_operand_inf = eq_1977 & eq_1978 | eq_1979 & eq_1980;
  assign and_reduce_2002 = &wide_exponent__2[7:0];
  assign has_pos_inf = ~(x_bexp__5 != MAX_EXPONENT__3 | ne_1983 | x_sign__1) | ~(y_bexp__5 != MAX_EXPONENT__4 | ne_1985 | y_sign__3);
  assign has_neg_inf = eq_1977 & eq_1978 & x_sign__1 | eq_1979 & eq_1980 & y_sign__3;
  assign fraction_shift__1 = rounding_carry ? fraction_shift__4 : fraction_shift__2;
  assign concat_2012 = {~(add_1895[25] | fraction_is_zero), add_1895[25], fraction_is_zero};
  assign shrl_2015 = rounded_fraction >> fraction_shift__1;
  assign is_result_nan = eq_1977 & ne_1983 | eq_1979 & ne_1985 | has_pos_inf & has_neg_inf;
  assign result_sign = x_sign__1 & y_sign__3 & concat_2012[0] | ~y_sign__3 & concat_2012[1] | y_sign__3 & concat_2012[2];
  assign result_fraction = shrl_2015[22:0];
  assign result_sign__1 = is_operand_inf ? ~has_pos_inf : result_sign;
  assign MAX_EXPONENT__2 = 8'hff;
  assign result_fraction__3 = result_fraction & {23{~(is_operand_inf | wide_exponent__2[8] | and_reduce_2002 | ~((|wide_exponent__2[8:1]) | wide_exponent__2[0]))}};
  assign FRACTION_HIGH_BIT = 23'h40_0000;
  assign result_sign__2 = ~is_result_nan & result_sign__1;
  assign result_exponent__2 = is_result_nan | is_operand_inf | wide_exponent__2[8] | and_reduce_2002 ? MAX_EXPONENT__2 : wide_exponent__2[7:0];
  assign result_fraction__4 = is_result_nan ? FRACTION_HIGH_BIT : result_fraction__3;
  assign out = {result_sign__2, result_exponent__2, result_fraction__4};
endmodule
