module COMP16 (x_a, x_b, wx);
  input  [15:0] x_a, x_b;
  output wx;
  wire [15:0] XOR;
  wire [7:0] temp;
  wire GT2_8,GT2_7,GT2_6,GT2_5,GT2_4,GT2_3,GT2_2,GT2_1;
  wire GT4_4,GT4_3,GT4_2,GT4_1;
  wire GT8_2,GT8_1;
  wire GT16_1;
  wire AND15_8,AND15_12,AND11_8,AND7_4; 
  
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[15]= x_a[15] ^ (!x_b[15]); //depth1
  assign XOR[14]= x_a[14] ^ (!x_b[14]);
  assign GT2_8 = (x_a[15] & (!x_b[15])) ^ (XOR[15] & x_a[14] & (!x_b[14]));//depth1
 
  assign XOR[13] = x_a[13] ^ (!x_b[13]);
  assign XOR[12] = x_a[12] ^ (!x_b[12]);
  assign GT2_7 = (x_a[13] & (!x_b[13])) ^ (XOR[13] & x_a[12] & (!x_b[12]));//depth1
  
  assign temp[4] = XOR[15] & XOR[14] & GT2_7;//depth2
  assign GT4_4 = temp[4] ^ GT2_8;//depth2
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[11]= x_a[11] ^ (!x_b[11]);
  assign XOR[10]= x_a[10] ^ (!x_b[10]);
  assign GT2_6 = (x_a[11] & (!x_b[11])) ^ (XOR[11] & x_a[10] & (!x_b[10]));//depth1
 
  assign XOR[9] = x_a[9] ^ (!x_b[9]);
  assign XOR[8] = x_a[8] ^ (!x_b[8]);
  assign GT2_5 = (x_a[9] & (!x_b[9])) ^ (XOR[9] & x_a[8] & (!x_b[8]));//depth1
  
  //assign temp[3] = XOR[11] & XOR[10] & GT2_5;//depth2
  //assign GT4_3 = temp[3] ^ GT2_6;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[6]= XOR[15] & XOR[14] & XOR[13] & XOR[12];//depth1
  assign AND15_12= (temp[6] & GT2_6) ^ (temp[6] & XOR[11] & XOR[10] & GT2_5);//depth2
  assign GT8_2 = AND15_12 ^ GT4_4;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[7]= x_a[7] ^ (!x_b[7]);
  assign XOR[6]= x_a[6] ^ (!x_b[6]);
  assign GT2_4 = (x_a[7] & (!x_b[7])) ^ (XOR[7] & x_a[6] & (!x_b[6]));//depth1
 
  assign XOR[5] = x_a[5] ^ (!x_b[5]);
  assign XOR[4] = x_a[4] ^ (!x_b[4]);
  assign GT2_3  = (x_a[5] & (!x_b[5])) ^ (XOR[5] & x_a[4] & (!x_b[4]));//depth1
  
  assign temp[2] = XOR[7] & XOR[6] & GT2_3;//depth2
  assign GT4_2 = temp[2] ^ GT2_4;//depth2
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[3]= x_a[3] ^ (!x_b[3]);
  assign XOR[2]= x_a[2] ^ (!x_b[2]);
  assign GT2_2 = (x_a[3] & (!x_b[3])) ^ (XOR[3] & x_a[2] & (!x_b[2]));//depth1
 
  assign XOR[1] = x_a[1] ^ (!x_b[1]);
  assign XOR[0] = x_a[0] ^ (!x_b[0]);
  assign GT2_1  = (x_a[1] & (!x_b[1])) ^ (XOR[1] & x_a[0] & (!x_b[0]));//depth1
  
  //assign temp[1] = XOR[3] & XOR[2] & GT2_1;//depth2
  //assign GT4_1 = temp[1] ^ GT2_2;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[5]= XOR[7] & XOR[6] & XOR[5] & XOR[4];//depth1
  assign AND7_4= (temp[5] & GT2_2) ^ (temp[5] & XOR[3] & XOR[2] & GT2_1);//depth2
  assign GT8_1 = AND7_4 ^ GT4_2;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign AND11_8= XOR[11] & XOR[10] & XOR[9] & XOR[8];//depth1
  assign temp[7]= AND11_8& temp[6];//depth2
  assign AND15_8=temp[7]&GT8_1;//depth3
  assign GT16_1 = AND15_8 ^ GT8_2;//depth3
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////


  assign wx = GT16_1;
endmodule



