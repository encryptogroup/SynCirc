module __f64sub__main(
  input wire [63:0] x,
  input wire [63:0] y,
  output wire [63:0] out
);
  wire [10:0] y_bexp__4;
  wire [10:0] x_bexp__4;
  wire [11:0] sum;
  wire [51:0] tuple_index_1850;
  wire [51:0] y_fraction__4;
  wire [10:0] y_bexp__5;
  wire [51:0] y_fraction__5;
  wire [10:0] incremented_sum__1;
  wire [56:0] wide_y;
  wire [10:0] x_bexpbs_difference__2;
  wire [10:0] x_bexp__5;
  wire [56:0] wide_y__1;
  wire [10:0] sub_1869;
  wire [51:0] x_fraction__1;
  wire [56:0] dropped;
  wire y_sign__2;
  wire [56:0] wide_x;
  wire tuple_index_1881;
  wire [56:0] wide_x__1;
  wire x_sign__1;
  wire y_sign__3;
  wire [56:0] neg_1887;
  wire [56:0] sticky;
  wire [56:0] xddend_y__1;
  wire [53:0] sel_1894;
  wire [54:0] add_1899;
  wire [56:0] concat_1902;
  wire [56:0] xbs_fraction__1;
  wire [56:0] reverse_1906;
  wire [57:0] one_hot_1907;
  wire [5:0] encode_1908;
  wire cancel__2;
  wire carry_bit;
  wire [56:0] leading_zeroes;
  wire [55:0] carry_fraction;
  wire [56:0] add_1925;
  wire [2:0] concat_1926;
  wire [55:0] carry_fraction__1;
  wire [55:0] cancel_fraction;
  wire [55:0] shifted_fraction;
  wire [2:0] normal_chunk;
  wire [2:0] fraction_shift__3;
  wire [1:0] half_way_chunk;
  wire [53:0] add_1941;
  wire do_round_up;
  wire [56:0] rounded_fraction;
  wire rounding_carry;
  wire [11:0] add_1952;
  wire [12:0] add_1960;
  wire [12:0] wide_exponent;
  wire [12:0] wide_exponent__1;
  wire [10:0] MAX_EXPONENT;
  wire [10:0] MAX_EXPONENT__1;
  wire [11:0] wide_exponent__2;
  wire [10:0] MAX_EXPONENT__3;
  wire [10:0] MAX_EXPONENT__4;
  wire eq_1981;
  wire eq_1982;
  wire eq_1983;
  wire eq_1984;
  wire ne_1987;
  wire ne_1989;
  wire fraction_is_zero;
  wire [2:0] fraction_shift__2;
  wire [2:0] fraction_shift__4;
  wire is_operand_inf;
  wire and_reduce_2006;
  wire has_pos_inf;
  wire has_neg_inf;
  wire [2:0] fraction_shift__1;
  wire [2:0] concat_2016;
  wire [56:0] shrl_2019;
  wire is_result_nan;
  wire result_sign;
  wire [51:0] result_fraction;
  wire result_sign__1;
  wire [10:0] MAX_EXPONENT__2;
  wire [51:0] result_fraction__3;
  wire [51:0] FRACTION_HIGH_BIT;
  wire result_sign__2;
  wire [10:0] result_exponent__2;
  wire [51:0] result_fraction__4;
  assign y_bexp__4 = y[62:52];
  assign x_bexp__4 = x[62:52];
  assign sum = {1'h0, x_bexp__4} + {1'h0, ~y_bexp__4};
  assign tuple_index_1850 = x[51:0];
  assign y_fraction__4 = y[51:0];
  assign y_bexp__5 = sum[11] ? y_bexp__4 : x_bexp__4;
  assign y_fraction__5 = sum[11] ? y_fraction__4 : tuple_index_1850;
  assign incremented_sum__1 = sum[10:0] + 11'h001;
  assign wide_y = {2'h1, y_fraction__5, 3'h0};
  assign x_bexpbs_difference__2 = sum[11] ? incremented_sum__1 : ~sum[10:0];
  assign x_bexp__5 = sum[11] ? x_bexp__4 : y_bexp__4;
  assign wide_y__1 = wide_y & {57{y_bexp__5 != 11'h000}};
  assign sub_1869 = 11'h039 - x_bexpbs_difference__2;
  assign x_fraction__1 = sum[11] ? tuple_index_1850 : y_fraction__4;
  assign dropped = sub_1869 >= 11'h039 ? 57'h000_0000_0000_0000 : wide_y__1 << sub_1869;
  assign y_sign__2 = y[63:63];
  assign wide_x = {2'h1, x_fraction__1, 3'h0};
  assign tuple_index_1881 = x[63:63];
  assign wide_x__1 = wide_x & {57{x_bexp__5 != 11'h000}};
  assign x_sign__1 = sum[11] ? tuple_index_1881 : ~y_sign__2;
  assign y_sign__3 = sum[11] ? ~y_sign__2 : tuple_index_1881;
  assign neg_1887 = -wide_x__1;
  assign sticky = {56'h00_0000_0000_0000, dropped[56:3] != 54'h00_0000_0000_0000};
  assign xddend_y__1 = (x_bexpbs_difference__2 >= 11'h039 ? 57'h000_0000_0000_0000 : wide_y__1 >> x_bexpbs_difference__2) | sticky;
  assign sel_1894 = x_sign__1 ^ y_sign__3 ? neg_1887[56:3] : wide_x__1[56:3];
  assign add_1899 = {{1{sel_1894[53]}}, sel_1894} + {1'h0, xddend_y__1[56:3]};
  assign concat_1902 = {add_1899[53:0], xddend_y__1[2:0]};
  assign xbs_fraction__1 = add_1899[54] ? -concat_1902 : concat_1902;
  assign reverse_1906 = {xbs_fraction__1[0], xbs_fraction__1[1], xbs_fraction__1[2], xbs_fraction__1[3], xbs_fraction__1[4], xbs_fraction__1[5], xbs_fraction__1[6], xbs_fraction__1[7], xbs_fraction__1[8], xbs_fraction__1[9], xbs_fraction__1[10], xbs_fraction__1[11], xbs_fraction__1[12], xbs_fraction__1[13], xbs_fraction__1[14], xbs_fraction__1[15], xbs_fraction__1[16], xbs_fraction__1[17], xbs_fraction__1[18], xbs_fraction__1[19], xbs_fraction__1[20], xbs_fraction__1[21], xbs_fraction__1[22], xbs_fraction__1[23], xbs_fraction__1[24], xbs_fraction__1[25], xbs_fraction__1[26], xbs_fraction__1[27], xbs_fraction__1[28], xbs_fraction__1[29], xbs_fraction__1[30], xbs_fraction__1[31], xbs_fraction__1[32], xbs_fraction__1[33], xbs_fraction__1[34], xbs_fraction__1[35], xbs_fraction__1[36], xbs_fraction__1[37], xbs_fraction__1[38], xbs_fraction__1[39], xbs_fraction__1[40], xbs_fraction__1[41], xbs_fraction__1[42], xbs_fraction__1[43], xbs_fraction__1[44], xbs_fraction__1[45], xbs_fraction__1[46], xbs_fraction__1[47], xbs_fraction__1[48], xbs_fraction__1[49], xbs_fraction__1[50], xbs_fraction__1[51], xbs_fraction__1[52], xbs_fraction__1[53], xbs_fraction__1[54], xbs_fraction__1[55], xbs_fraction__1[56]};
  assign one_hot_1907 = {reverse_1906[56:0] == 57'h000_0000_0000_0000, reverse_1906[56] && reverse_1906[55:0] == 56'h00_0000_0000_0000, reverse_1906[55] && reverse_1906[54:0] == 55'h00_0000_0000_0000, reverse_1906[54] && reverse_1906[53:0] == 54'h00_0000_0000_0000, reverse_1906[53] && reverse_1906[52:0] == 53'h00_0000_0000_0000, reverse_1906[52] && reverse_1906[51:0] == 52'h0_0000_0000_0000, reverse_1906[51] && reverse_1906[50:0] == 51'h0_0000_0000_0000, reverse_1906[50] && reverse_1906[49:0] == 50'h0_0000_0000_0000, reverse_1906[49] && reverse_1906[48:0] == 49'h0_0000_0000_0000, reverse_1906[48] && reverse_1906[47:0] == 48'h0000_0000_0000, reverse_1906[47] && reverse_1906[46:0] == 47'h0000_0000_0000, reverse_1906[46] && reverse_1906[45:0] == 46'h0000_0000_0000, reverse_1906[45] && reverse_1906[44:0] == 45'h0000_0000_0000, reverse_1906[44] && reverse_1906[43:0] == 44'h000_0000_0000, reverse_1906[43] && reverse_1906[42:0] == 43'h000_0000_0000, reverse_1906[42] && reverse_1906[41:0] == 42'h000_0000_0000, reverse_1906[41] && reverse_1906[40:0] == 41'h000_0000_0000, reverse_1906[40] && reverse_1906[39:0] == 40'h00_0000_0000, reverse_1906[39] && reverse_1906[38:0] == 39'h00_0000_0000, reverse_1906[38] && reverse_1906[37:0] == 38'h00_0000_0000, reverse_1906[37] && reverse_1906[36:0] == 37'h00_0000_0000, reverse_1906[36] && reverse_1906[35:0] == 36'h0_0000_0000, reverse_1906[35] && reverse_1906[34:0] == 35'h0_0000_0000, reverse_1906[34] && reverse_1906[33:0] == 34'h0_0000_0000, reverse_1906[33] && reverse_1906[32:0] == 33'h0_0000_0000, reverse_1906[32] && reverse_1906[31:0] == 32'h0000_0000, reverse_1906[31] && reverse_1906[30:0] == 31'h0000_0000, reverse_1906[30] && reverse_1906[29:0] == 30'h0000_0000, reverse_1906[29] && reverse_1906[28:0] == 29'h0000_0000, reverse_1906[28] && reverse_1906[27:0] == 28'h000_0000, reverse_1906[27] && reverse_1906[26:0] == 27'h000_0000, reverse_1906[26] && reverse_1906[25:0] == 26'h000_0000, reverse_1906[25] && reverse_1906[24:0] == 25'h000_0000, reverse_1906[24] && reverse_1906[23:0] == 24'h00_0000, reverse_1906[23] && reverse_1906[22:0] == 23'h00_0000, reverse_1906[22] && reverse_1906[21:0] == 22'h00_0000, reverse_1906[21] && reverse_1906[20:0] == 21'h00_0000, reverse_1906[20] && reverse_1906[19:0] == 20'h0_0000, reverse_1906[19] && reverse_1906[18:0] == 19'h0_0000, reverse_1906[18] && reverse_1906[17:0] == 18'h0_0000, reverse_1906[17] && reverse_1906[16:0] == 17'h0_0000, reverse_1906[16] && reverse_1906[15:0] == 16'h0000, reverse_1906[15] && reverse_1906[14:0] == 15'h0000, reverse_1906[14] && reverse_1906[13:0] == 14'h0000, reverse_1906[13] && reverse_1906[12:0] == 13'h0000, reverse_1906[12] && reverse_1906[11:0] == 12'h000, reverse_1906[11] && reverse_1906[10:0] == 11'h000, reverse_1906[10] && reverse_1906[9:0] == 10'h000, reverse_1906[9] && reverse_1906[8:0] == 9'h000, reverse_1906[8] && reverse_1906[7:0] == 8'h00, reverse_1906[7] && reverse_1906[6:0] == 7'h00, reverse_1906[6] && reverse_1906[5:0] == 6'h00, reverse_1906[5] && reverse_1906[4:0] == 5'h00, reverse_1906[4] && reverse_1906[3:0] == 4'h0, reverse_1906[3] && reverse_1906[2:0] == 3'h0, reverse_1906[2] && reverse_1906[1:0] == 2'h0, reverse_1906[1] && !reverse_1906[0], reverse_1906[0]};
  assign encode_1908 = {one_hot_1907[32] | one_hot_1907[33] | one_hot_1907[34] | one_hot_1907[35] | one_hot_1907[36] | one_hot_1907[37] | one_hot_1907[38] | one_hot_1907[39] | one_hot_1907[40] | one_hot_1907[41] | one_hot_1907[42] | one_hot_1907[43] | one_hot_1907[44] | one_hot_1907[45] | one_hot_1907[46] | one_hot_1907[47] | one_hot_1907[48] | one_hot_1907[49] | one_hot_1907[50] | one_hot_1907[51] | one_hot_1907[52] | one_hot_1907[53] | one_hot_1907[54] | one_hot_1907[55] | one_hot_1907[56] | one_hot_1907[57], one_hot_1907[16] | one_hot_1907[17] | one_hot_1907[18] | one_hot_1907[19] | one_hot_1907[20] | one_hot_1907[21] | one_hot_1907[22] | one_hot_1907[23] | one_hot_1907[24] | one_hot_1907[25] | one_hot_1907[26] | one_hot_1907[27] | one_hot_1907[28] | one_hot_1907[29] | one_hot_1907[30] | one_hot_1907[31] | one_hot_1907[48] | one_hot_1907[49] | one_hot_1907[50] | one_hot_1907[51] | one_hot_1907[52] | one_hot_1907[53] | one_hot_1907[54] | one_hot_1907[55] | one_hot_1907[56] | one_hot_1907[57], one_hot_1907[8] | one_hot_1907[9] | one_hot_1907[10] | one_hot_1907[11] | one_hot_1907[12] | one_hot_1907[13] | one_hot_1907[14] | one_hot_1907[15] | one_hot_1907[24] | one_hot_1907[25] | one_hot_1907[26] | one_hot_1907[27] | one_hot_1907[28] | one_hot_1907[29] | one_hot_1907[30] | one_hot_1907[31] | one_hot_1907[40] | one_hot_1907[41] | one_hot_1907[42] | one_hot_1907[43] | one_hot_1907[44] | one_hot_1907[45] | one_hot_1907[46] | one_hot_1907[47] | one_hot_1907[56] | one_hot_1907[57], one_hot_1907[4] | one_hot_1907[5] | one_hot_1907[6] | one_hot_1907[7] | one_hot_1907[12] | one_hot_1907[13] | one_hot_1907[14] | one_hot_1907[15] | one_hot_1907[20] | one_hot_1907[21] | one_hot_1907[22] | one_hot_1907[23] | one_hot_1907[28] | one_hot_1907[29] | one_hot_1907[30] | one_hot_1907[31] | one_hot_1907[36] | one_hot_1907[37] | one_hot_1907[38] | one_hot_1907[39] | one_hot_1907[44] | one_hot_1907[45] | one_hot_1907[46] | one_hot_1907[47] | one_hot_1907[52] | one_hot_1907[53] | one_hot_1907[54] | one_hot_1907[55], one_hot_1907[2] | one_hot_1907[3] | one_hot_1907[6] | one_hot_1907[7] | one_hot_1907[10] | one_hot_1907[11] | one_hot_1907[14] | one_hot_1907[15] | one_hot_1907[18] | one_hot_1907[19] | one_hot_1907[22] | one_hot_1907[23] | one_hot_1907[26] | one_hot_1907[27] | one_hot_1907[30] | one_hot_1907[31] | one_hot_1907[34] | one_hot_1907[35] | one_hot_1907[38] | one_hot_1907[39] | one_hot_1907[42] | one_hot_1907[43] | one_hot_1907[46] | one_hot_1907[47] | one_hot_1907[50] | one_hot_1907[51] | one_hot_1907[54] | one_hot_1907[55], one_hot_1907[1] | one_hot_1907[3] | one_hot_1907[5] | one_hot_1907[7] | one_hot_1907[9] | one_hot_1907[11] | one_hot_1907[13] | one_hot_1907[15] | one_hot_1907[17] | one_hot_1907[19] | one_hot_1907[21] | one_hot_1907[23] | one_hot_1907[25] | one_hot_1907[27] | one_hot_1907[29] | one_hot_1907[31] | one_hot_1907[33] | one_hot_1907[35] | one_hot_1907[37] | one_hot_1907[39] | one_hot_1907[41] | one_hot_1907[43] | one_hot_1907[45] | one_hot_1907[47] | one_hot_1907[49] | one_hot_1907[51] | one_hot_1907[53] | one_hot_1907[55] | one_hot_1907[57]};
  assign cancel__2 = |encode_1908[5:1];
  assign carry_bit = xbs_fraction__1[56];
  assign leading_zeroes = {51'h0_0000_0000_0000, encode_1908};
  assign carry_fraction = xbs_fraction__1[56:1];
  assign add_1925 = leading_zeroes + 57'h1ff_ffff_ffff_ffff;
  assign concat_1926 = {~(carry_bit | cancel__2), ~(carry_bit | ~cancel__2), ~(~carry_bit | cancel__2)};
  assign carry_fraction__1 = carry_fraction | {55'h00_0000_0000_0000, xbs_fraction__1[0]};
  assign cancel_fraction = add_1925 >= 57'h000_0000_0000_0038 ? 56'h00_0000_0000_0000 : xbs_fraction__1[55:0] << add_1925;
  assign shifted_fraction = carry_fraction__1 & {56{concat_1926[0]}} | cancel_fraction & {56{concat_1926[1]}} | xbs_fraction__1[55:0] & {56{concat_1926[2]}};
  assign normal_chunk = shifted_fraction[2:0];
  assign fraction_shift__3 = 3'h4;
  assign half_way_chunk = shifted_fraction[3:2];
  assign add_1941 = {1'h0, shifted_fraction[55:3]} + 54'h00_0000_0000_0001;
  assign do_round_up = normal_chunk > fraction_shift__3 | half_way_chunk == 2'h3;
  assign rounded_fraction = do_round_up ? {add_1941, normal_chunk} : {1'h0, shifted_fraction};
  assign rounding_carry = rounded_fraction[56];
  assign add_1952 = {1'h0, x_bexp__5} + {11'h000, rounding_carry};
  assign add_1960 = {1'h0, add_1952} + 13'h0001;
  assign wide_exponent = add_1960 - {7'h00, encode_1908};
  assign wide_exponent__1 = wide_exponent & {13{add_1899 != 55'h00_0000_0000_0000 | xddend_y__1[2:0] != 3'h0}};
  assign MAX_EXPONENT = 11'h7ff;
  assign MAX_EXPONENT__1 = 11'h7ff;
  assign wide_exponent__2 = wide_exponent__1[11:0] & {12{~wide_exponent__1[12]}};
  assign MAX_EXPONENT__3 = 11'h7ff;
  assign MAX_EXPONENT__4 = 11'h7ff;
  assign eq_1981 = x_bexp__5 == MAX_EXPONENT;
  assign eq_1982 = x_fraction__1 == 52'h0_0000_0000_0000;
  assign eq_1983 = y_bexp__5 == MAX_EXPONENT__1;
  assign eq_1984 = y_fraction__5 == 52'h0_0000_0000_0000;
  assign ne_1987 = x_fraction__1 != 52'h0_0000_0000_0000;
  assign ne_1989 = y_fraction__5 != 52'h0_0000_0000_0000;
  assign fraction_is_zero = add_1899 == 55'h00_0000_0000_0000 & xddend_y__1[2:0] == 3'h0;
  assign fraction_shift__2 = 3'h3;
  assign fraction_shift__4 = 3'h4;
  assign is_operand_inf = eq_1981 & eq_1982 | eq_1983 & eq_1984;
  assign and_reduce_2006 = &wide_exponent__2[10:0];
  assign has_pos_inf = ~(x_bexp__5 != MAX_EXPONENT__3 | ne_1987 | x_sign__1) | ~(y_bexp__5 != MAX_EXPONENT__4 | ne_1989 | y_sign__3);
  assign has_neg_inf = eq_1981 & eq_1982 & x_sign__1 | eq_1983 & eq_1984 & y_sign__3;
  assign fraction_shift__1 = rounding_carry ? fraction_shift__4 : fraction_shift__2;
  assign concat_2016 = {~(add_1899[54] | fraction_is_zero), add_1899[54], fraction_is_zero};
  assign shrl_2019 = rounded_fraction >> fraction_shift__1;
  assign is_result_nan = eq_1981 & ne_1987 | eq_1983 & ne_1989 | has_pos_inf & has_neg_inf;
  assign result_sign = x_sign__1 & y_sign__3 & concat_2016[0] | ~y_sign__3 & concat_2016[1] | y_sign__3 & concat_2016[2];
  assign result_fraction = shrl_2019[51:0];
  assign result_sign__1 = is_operand_inf ? ~has_pos_inf : result_sign;
  assign MAX_EXPONENT__2 = 11'h7ff;
  assign result_fraction__3 = result_fraction & {52{~(is_operand_inf | wide_exponent__2[11] | and_reduce_2006 | ~((|wide_exponent__2[11:1]) | wide_exponent__2[0]))}};
  assign FRACTION_HIGH_BIT = 52'h8_0000_0000_0000;
  assign result_sign__2 = ~is_result_nan & result_sign__1;
  assign result_exponent__2 = is_result_nan | is_operand_inf | wide_exponent__2[11] | and_reduce_2006 ? MAX_EXPONENT__2 : wide_exponent__2[10:0];
  assign result_fraction__4 = is_result_nan ? FRACTION_HIGH_BIT : result_fraction__3;
  assign out = {result_sign__2, result_exponent__2, result_fraction__4};
endmodule
