module main(input [31:0] a, input [31:0] b, output [31:0] y);
   f32add f32add(a, b, y);
endmodule // main
