module __f64add__main(
  input wire [63:0] x,
  input wire [63:0] y,
  output wire [63:0] out
);
  wire [10:0] y_bexp__1;
  wire [10:0] x_bexp__1;
  wire [11:0] sum;
  wire [51:0] tuple_index_1624;
  wire [51:0] tuple_index_1625;
  wire [10:0] y_bexp__2;
  wire [51:0] y_fraction__1;
  wire [10:0] incremented_sum__1;
  wire [56:0] wide_y;
  wire [10:0] x_bexpbs_difference__1;
  wire [10:0] x_bexp__2;
  wire [56:0] wide_y__1;
  wire [10:0] sub_1643;
  wire [51:0] x_fraction__2;
  wire [56:0] dropped;
  wire [56:0] wide_x;
  wire tuple_index_1653;
  wire tuple_index_1654;
  wire [56:0] wide_x__1;
  wire x_sign__2;
  wire y_sign__2;
  wire [56:0] neg_1660;
  wire [56:0] sticky;
  wire [56:0] xddend_y__2;
  wire [53:0] sel_1667;
  wire [54:0] add_1672;
  wire [56:0] concat_1675;
  wire [56:0] xbs_fraction__2;
  wire [56:0] reverse_1679;
  wire [57:0] one_hot_1680;
  wire [5:0] encode_1681;
  wire cancel__2;
  wire carry_bit;
  wire [56:0] leading_zeroes;
  wire [55:0] carry_fraction;
  wire [56:0] add_1698;
  wire [2:0] concat_1699;
  wire [55:0] carry_fraction__1;
  wire [55:0] cancel_fraction;
  wire [55:0] shifted_fraction;
  wire [2:0] normal_chunk;
  wire [2:0] fraction_shift__3;
  wire [1:0] half_way_chunk;
  wire [53:0] add_1714;
  wire do_round_up;
  wire [56:0] rounded_fraction;
  wire rounding_carry;
  wire [11:0] add_1725;
  wire [12:0] add_1733;
  wire [12:0] wide_exponent;
  wire [12:0] wide_exponent__1;
  wire [10:0] MAX_EXPONENT;
  wire [10:0] MAX_EXPONENT__1;
  wire [11:0] wide_exponent__2;
  wire [10:0] MAX_EXPONENT__3;
  wire [10:0] MAX_EXPONENT__4;
  wire eq_1754;
  wire eq_1755;
  wire eq_1756;
  wire eq_1757;
  wire ne_1760;
  wire ne_1762;
  wire fraction_is_zero;
  wire [2:0] fraction_shift__2;
  wire [2:0] fraction_shift__4;
  wire is_operand_inf;
  wire and_reduce_1779;
  wire has_pos_inf;
  wire has_neg_inf;
  wire [2:0] fraction_shift__1;
  wire [2:0] concat_1789;
  wire [56:0] shrl_1792;
  wire is_result_nan;
  wire result_sign;
  wire [51:0] result_fraction;
  wire result_sign__1;
  wire [10:0] MAX_EXPONENT__2;
  wire [51:0] result_fraction__3;
  wire [51:0] FRACTION_HIGH_BIT;
  wire result_sign__2;
  wire [10:0] result_exponent__2;
  wire [51:0] result_fraction__4;
  assign y_bexp__1 = y[62:52];
  assign x_bexp__1 = x[62:52];
  assign sum = {1'h0, x_bexp__1} + {1'h0, ~y_bexp__1};
  assign tuple_index_1624 = x[51:0];
  assign tuple_index_1625 = y[51:0];
  assign y_bexp__2 = sum[11] ? y_bexp__1 : x_bexp__1;
  assign y_fraction__1 = sum[11] ? tuple_index_1625 : tuple_index_1624;
  assign incremented_sum__1 = sum[10:0] + 11'h001;
  assign wide_y = {2'h1, y_fraction__1, 3'h0};
  assign x_bexpbs_difference__1 = sum[11] ? incremented_sum__1 : ~sum[10:0];
  assign x_bexp__2 = sum[11] ? x_bexp__1 : y_bexp__1;
  assign wide_y__1 = wide_y & {57{y_bexp__2 != 11'h000}};
  assign sub_1643 = 11'h039 - x_bexpbs_difference__1;
  assign x_fraction__2 = sum[11] ? tuple_index_1624 : tuple_index_1625;
  assign dropped = sub_1643 >= 11'h039 ? 57'h000_0000_0000_0000 : wide_y__1 << sub_1643;
  assign wide_x = {2'h1, x_fraction__2, 3'h0};
  assign tuple_index_1653 = y[63:63];
  assign tuple_index_1654 = x[63:63];
  assign wide_x__1 = wide_x & {57{x_bexp__2 != 11'h000}};
  assign x_sign__2 = sum[11] ? tuple_index_1654 : tuple_index_1653;
  assign y_sign__2 = sum[11] ? tuple_index_1653 : tuple_index_1654;
  assign neg_1660 = -wide_x__1;
  assign sticky = {56'h00_0000_0000_0000, dropped[56:3] != 54'h00_0000_0000_0000};
  assign xddend_y__2 = (x_bexpbs_difference__1 >= 11'h039 ? 57'h000_0000_0000_0000 : wide_y__1 >> x_bexpbs_difference__1) | sticky;
  assign sel_1667 = x_sign__2 ^ y_sign__2 ? neg_1660[56:3] : wide_x__1[56:3];
  assign add_1672 = {{1{sel_1667[53]}}, sel_1667} + {1'h0, xddend_y__2[56:3]};
  assign concat_1675 = {add_1672[53:0], xddend_y__2[2:0]};
  assign xbs_fraction__2 = add_1672[54] ? -concat_1675 : concat_1675;
  assign reverse_1679 = {xbs_fraction__2[0], xbs_fraction__2[1], xbs_fraction__2[2], xbs_fraction__2[3], xbs_fraction__2[4], xbs_fraction__2[5], xbs_fraction__2[6], xbs_fraction__2[7], xbs_fraction__2[8], xbs_fraction__2[9], xbs_fraction__2[10], xbs_fraction__2[11], xbs_fraction__2[12], xbs_fraction__2[13], xbs_fraction__2[14], xbs_fraction__2[15], xbs_fraction__2[16], xbs_fraction__2[17], xbs_fraction__2[18], xbs_fraction__2[19], xbs_fraction__2[20], xbs_fraction__2[21], xbs_fraction__2[22], xbs_fraction__2[23], xbs_fraction__2[24], xbs_fraction__2[25], xbs_fraction__2[26], xbs_fraction__2[27], xbs_fraction__2[28], xbs_fraction__2[29], xbs_fraction__2[30], xbs_fraction__2[31], xbs_fraction__2[32], xbs_fraction__2[33], xbs_fraction__2[34], xbs_fraction__2[35], xbs_fraction__2[36], xbs_fraction__2[37], xbs_fraction__2[38], xbs_fraction__2[39], xbs_fraction__2[40], xbs_fraction__2[41], xbs_fraction__2[42], xbs_fraction__2[43], xbs_fraction__2[44], xbs_fraction__2[45], xbs_fraction__2[46], xbs_fraction__2[47], xbs_fraction__2[48], xbs_fraction__2[49], xbs_fraction__2[50], xbs_fraction__2[51], xbs_fraction__2[52], xbs_fraction__2[53], xbs_fraction__2[54], xbs_fraction__2[55], xbs_fraction__2[56]};
  assign one_hot_1680 = {reverse_1679[56:0] == 57'h000_0000_0000_0000, reverse_1679[56] && reverse_1679[55:0] == 56'h00_0000_0000_0000, reverse_1679[55] && reverse_1679[54:0] == 55'h00_0000_0000_0000, reverse_1679[54] && reverse_1679[53:0] == 54'h00_0000_0000_0000, reverse_1679[53] && reverse_1679[52:0] == 53'h00_0000_0000_0000, reverse_1679[52] && reverse_1679[51:0] == 52'h0_0000_0000_0000, reverse_1679[51] && reverse_1679[50:0] == 51'h0_0000_0000_0000, reverse_1679[50] && reverse_1679[49:0] == 50'h0_0000_0000_0000, reverse_1679[49] && reverse_1679[48:0] == 49'h0_0000_0000_0000, reverse_1679[48] && reverse_1679[47:0] == 48'h0000_0000_0000, reverse_1679[47] && reverse_1679[46:0] == 47'h0000_0000_0000, reverse_1679[46] && reverse_1679[45:0] == 46'h0000_0000_0000, reverse_1679[45] && reverse_1679[44:0] == 45'h0000_0000_0000, reverse_1679[44] && reverse_1679[43:0] == 44'h000_0000_0000, reverse_1679[43] && reverse_1679[42:0] == 43'h000_0000_0000, reverse_1679[42] && reverse_1679[41:0] == 42'h000_0000_0000, reverse_1679[41] && reverse_1679[40:0] == 41'h000_0000_0000, reverse_1679[40] && reverse_1679[39:0] == 40'h00_0000_0000, reverse_1679[39] && reverse_1679[38:0] == 39'h00_0000_0000, reverse_1679[38] && reverse_1679[37:0] == 38'h00_0000_0000, reverse_1679[37] && reverse_1679[36:0] == 37'h00_0000_0000, reverse_1679[36] && reverse_1679[35:0] == 36'h0_0000_0000, reverse_1679[35] && reverse_1679[34:0] == 35'h0_0000_0000, reverse_1679[34] && reverse_1679[33:0] == 34'h0_0000_0000, reverse_1679[33] && reverse_1679[32:0] == 33'h0_0000_0000, reverse_1679[32] && reverse_1679[31:0] == 32'h0000_0000, reverse_1679[31] && reverse_1679[30:0] == 31'h0000_0000, reverse_1679[30] && reverse_1679[29:0] == 30'h0000_0000, reverse_1679[29] && reverse_1679[28:0] == 29'h0000_0000, reverse_1679[28] && reverse_1679[27:0] == 28'h000_0000, reverse_1679[27] && reverse_1679[26:0] == 27'h000_0000, reverse_1679[26] && reverse_1679[25:0] == 26'h000_0000, reverse_1679[25] && reverse_1679[24:0] == 25'h000_0000, reverse_1679[24] && reverse_1679[23:0] == 24'h00_0000, reverse_1679[23] && reverse_1679[22:0] == 23'h00_0000, reverse_1679[22] && reverse_1679[21:0] == 22'h00_0000, reverse_1679[21] && reverse_1679[20:0] == 21'h00_0000, reverse_1679[20] && reverse_1679[19:0] == 20'h0_0000, reverse_1679[19] && reverse_1679[18:0] == 19'h0_0000, reverse_1679[18] && reverse_1679[17:0] == 18'h0_0000, reverse_1679[17] && reverse_1679[16:0] == 17'h0_0000, reverse_1679[16] && reverse_1679[15:0] == 16'h0000, reverse_1679[15] && reverse_1679[14:0] == 15'h0000, reverse_1679[14] && reverse_1679[13:0] == 14'h0000, reverse_1679[13] && reverse_1679[12:0] == 13'h0000, reverse_1679[12] && reverse_1679[11:0] == 12'h000, reverse_1679[11] && reverse_1679[10:0] == 11'h000, reverse_1679[10] && reverse_1679[9:0] == 10'h000, reverse_1679[9] && reverse_1679[8:0] == 9'h000, reverse_1679[8] && reverse_1679[7:0] == 8'h00, reverse_1679[7] && reverse_1679[6:0] == 7'h00, reverse_1679[6] && reverse_1679[5:0] == 6'h00, reverse_1679[5] && reverse_1679[4:0] == 5'h00, reverse_1679[4] && reverse_1679[3:0] == 4'h0, reverse_1679[3] && reverse_1679[2:0] == 3'h0, reverse_1679[2] && reverse_1679[1:0] == 2'h0, reverse_1679[1] && !reverse_1679[0], reverse_1679[0]};
  assign encode_1681 = {one_hot_1680[32] | one_hot_1680[33] | one_hot_1680[34] | one_hot_1680[35] | one_hot_1680[36] | one_hot_1680[37] | one_hot_1680[38] | one_hot_1680[39] | one_hot_1680[40] | one_hot_1680[41] | one_hot_1680[42] | one_hot_1680[43] | one_hot_1680[44] | one_hot_1680[45] | one_hot_1680[46] | one_hot_1680[47] | one_hot_1680[48] | one_hot_1680[49] | one_hot_1680[50] | one_hot_1680[51] | one_hot_1680[52] | one_hot_1680[53] | one_hot_1680[54] | one_hot_1680[55] | one_hot_1680[56] | one_hot_1680[57], one_hot_1680[16] | one_hot_1680[17] | one_hot_1680[18] | one_hot_1680[19] | one_hot_1680[20] | one_hot_1680[21] | one_hot_1680[22] | one_hot_1680[23] | one_hot_1680[24] | one_hot_1680[25] | one_hot_1680[26] | one_hot_1680[27] | one_hot_1680[28] | one_hot_1680[29] | one_hot_1680[30] | one_hot_1680[31] | one_hot_1680[48] | one_hot_1680[49] | one_hot_1680[50] | one_hot_1680[51] | one_hot_1680[52] | one_hot_1680[53] | one_hot_1680[54] | one_hot_1680[55] | one_hot_1680[56] | one_hot_1680[57], one_hot_1680[8] | one_hot_1680[9] | one_hot_1680[10] | one_hot_1680[11] | one_hot_1680[12] | one_hot_1680[13] | one_hot_1680[14] | one_hot_1680[15] | one_hot_1680[24] | one_hot_1680[25] | one_hot_1680[26] | one_hot_1680[27] | one_hot_1680[28] | one_hot_1680[29] | one_hot_1680[30] | one_hot_1680[31] | one_hot_1680[40] | one_hot_1680[41] | one_hot_1680[42] | one_hot_1680[43] | one_hot_1680[44] | one_hot_1680[45] | one_hot_1680[46] | one_hot_1680[47] | one_hot_1680[56] | one_hot_1680[57], one_hot_1680[4] | one_hot_1680[5] | one_hot_1680[6] | one_hot_1680[7] | one_hot_1680[12] | one_hot_1680[13] | one_hot_1680[14] | one_hot_1680[15] | one_hot_1680[20] | one_hot_1680[21] | one_hot_1680[22] | one_hot_1680[23] | one_hot_1680[28] | one_hot_1680[29] | one_hot_1680[30] | one_hot_1680[31] | one_hot_1680[36] | one_hot_1680[37] | one_hot_1680[38] | one_hot_1680[39] | one_hot_1680[44] | one_hot_1680[45] | one_hot_1680[46] | one_hot_1680[47] | one_hot_1680[52] | one_hot_1680[53] | one_hot_1680[54] | one_hot_1680[55], one_hot_1680[2] | one_hot_1680[3] | one_hot_1680[6] | one_hot_1680[7] | one_hot_1680[10] | one_hot_1680[11] | one_hot_1680[14] | one_hot_1680[15] | one_hot_1680[18] | one_hot_1680[19] | one_hot_1680[22] | one_hot_1680[23] | one_hot_1680[26] | one_hot_1680[27] | one_hot_1680[30] | one_hot_1680[31] | one_hot_1680[34] | one_hot_1680[35] | one_hot_1680[38] | one_hot_1680[39] | one_hot_1680[42] | one_hot_1680[43] | one_hot_1680[46] | one_hot_1680[47] | one_hot_1680[50] | one_hot_1680[51] | one_hot_1680[54] | one_hot_1680[55], one_hot_1680[1] | one_hot_1680[3] | one_hot_1680[5] | one_hot_1680[7] | one_hot_1680[9] | one_hot_1680[11] | one_hot_1680[13] | one_hot_1680[15] | one_hot_1680[17] | one_hot_1680[19] | one_hot_1680[21] | one_hot_1680[23] | one_hot_1680[25] | one_hot_1680[27] | one_hot_1680[29] | one_hot_1680[31] | one_hot_1680[33] | one_hot_1680[35] | one_hot_1680[37] | one_hot_1680[39] | one_hot_1680[41] | one_hot_1680[43] | one_hot_1680[45] | one_hot_1680[47] | one_hot_1680[49] | one_hot_1680[51] | one_hot_1680[53] | one_hot_1680[55] | one_hot_1680[57]};
  assign cancel__2 = |encode_1681[5:1];
  assign carry_bit = xbs_fraction__2[56];
  assign leading_zeroes = {51'h0_0000_0000_0000, encode_1681};
  assign carry_fraction = xbs_fraction__2[56:1];
  assign add_1698 = leading_zeroes + 57'h1ff_ffff_ffff_ffff;
  assign concat_1699 = {~(carry_bit | cancel__2), ~(carry_bit | ~cancel__2), ~(~carry_bit | cancel__2)};
  assign carry_fraction__1 = carry_fraction | {55'h00_0000_0000_0000, xbs_fraction__2[0]};
  assign cancel_fraction = add_1698 >= 57'h000_0000_0000_0038 ? 56'h00_0000_0000_0000 : xbs_fraction__2[55:0] << add_1698;
  assign shifted_fraction = carry_fraction__1 & {56{concat_1699[0]}} | cancel_fraction & {56{concat_1699[1]}} | xbs_fraction__2[55:0] & {56{concat_1699[2]}};
  assign normal_chunk = shifted_fraction[2:0];
  assign fraction_shift__3 = 3'h4;
  assign half_way_chunk = shifted_fraction[3:2];
  assign add_1714 = {1'h0, shifted_fraction[55:3]} + 54'h00_0000_0000_0001;
  assign do_round_up = normal_chunk > fraction_shift__3 | half_way_chunk == 2'h3;
  assign rounded_fraction = do_round_up ? {add_1714, normal_chunk} : {1'h0, shifted_fraction};
  assign rounding_carry = rounded_fraction[56];
  assign add_1725 = {1'h0, x_bexp__2} + {11'h000, rounding_carry};
  assign add_1733 = {1'h0, add_1725} + 13'h0001;
  assign wide_exponent = add_1733 - {7'h00, encode_1681};
  assign wide_exponent__1 = wide_exponent & {13{add_1672 != 55'h00_0000_0000_0000 | xddend_y__2[2:0] != 3'h0}};
  assign MAX_EXPONENT = 11'h7ff;
  assign MAX_EXPONENT__1 = 11'h7ff;
  assign wide_exponent__2 = wide_exponent__1[11:0] & {12{~wide_exponent__1[12]}};
  assign MAX_EXPONENT__3 = 11'h7ff;
  assign MAX_EXPONENT__4 = 11'h7ff;
  assign eq_1754 = x_bexp__2 == MAX_EXPONENT;
  assign eq_1755 = x_fraction__2 == 52'h0_0000_0000_0000;
  assign eq_1756 = y_bexp__2 == MAX_EXPONENT__1;
  assign eq_1757 = y_fraction__1 == 52'h0_0000_0000_0000;
  assign ne_1760 = x_fraction__2 != 52'h0_0000_0000_0000;
  assign ne_1762 = y_fraction__1 != 52'h0_0000_0000_0000;
  assign fraction_is_zero = add_1672 == 55'h00_0000_0000_0000 & xddend_y__2[2:0] == 3'h0;
  assign fraction_shift__2 = 3'h3;
  assign fraction_shift__4 = 3'h4;
  assign is_operand_inf = eq_1754 & eq_1755 | eq_1756 & eq_1757;
  assign and_reduce_1779 = &wide_exponent__2[10:0];
  assign has_pos_inf = ~(x_bexp__2 != MAX_EXPONENT__3 | ne_1760 | x_sign__2) | ~(y_bexp__2 != MAX_EXPONENT__4 | ne_1762 | y_sign__2);
  assign has_neg_inf = eq_1754 & eq_1755 & x_sign__2 | eq_1756 & eq_1757 & y_sign__2;
  assign fraction_shift__1 = rounding_carry ? fraction_shift__4 : fraction_shift__2;
  assign concat_1789 = {~(add_1672[54] | fraction_is_zero), add_1672[54], fraction_is_zero};
  assign shrl_1792 = rounded_fraction >> fraction_shift__1;
  assign is_result_nan = eq_1754 & ne_1760 | eq_1756 & ne_1762 | has_pos_inf & has_neg_inf;
  assign result_sign = x_sign__2 & y_sign__2 & concat_1789[0] | ~y_sign__2 & concat_1789[1] | y_sign__2 & concat_1789[2];
  assign result_fraction = shrl_1792[51:0];
  assign result_sign__1 = is_operand_inf ? ~has_pos_inf : result_sign;
  assign MAX_EXPONENT__2 = 11'h7ff;
  assign result_fraction__3 = result_fraction & {52{~(is_operand_inf | wide_exponent__2[11] | and_reduce_1779 | ~((|wide_exponent__2[11:1]) | wide_exponent__2[0]))}};
  assign FRACTION_HIGH_BIT = 52'h8_0000_0000_0000;
  assign result_sign__2 = ~is_result_nan & result_sign__1;
  assign result_exponent__2 = is_result_nan | is_operand_inf | wide_exponent__2[11] | and_reduce_1779 ? MAX_EXPONENT__2 : wide_exponent__2[10:0];
  assign result_fraction__4 = is_result_nan ? FRACTION_HIGH_BIT : result_fraction__3;
  assign out = {result_sign__2, result_exponent__2, result_fraction__4};
endmodule
