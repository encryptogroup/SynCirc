module main(input [31:0] a, input [31:0] b, output [31:0] y);
   f32mul f32mul(a, b, y);
endmodule // main
