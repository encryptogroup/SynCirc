module COMP32 (x_a, x_b, wx);
  input  [31:0] x_a, x_b;
  output wx;
  wire [31:0] XOR;
  wire [15:0] temp;
  wire GT2_16,GT2_15,GT2_14,GT2_13,GT2_12,GT2_11,GT2_10,GT2_9,GT2_8,GT2_7,GT2_6,GT2_5,GT2_4,GT2_3,GT2_2,GT2_1;
  wire GT4_8,GT4_7,GT4_6,GT4_5,GT4_4,GT4_3,GT4_2,GT4_1;
  wire GT8_4,GT8_3,GT8_2,GT8_1;
  wire GT16_2,GT16_1;
  wire GT32_1;
  wire AND31_28,AND23_20,AND15_12,AND19_16,AND27_24,AND31_16,AND11_8,AND7_4,AND31_24; 
  
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[31]= x_a[31] ^ (!x_b[31]);
  assign XOR[30]= x_a[30] ^ (!x_b[30]);
  assign GT2_16 = (x_a[31] & (!x_b[31])) ^ (XOR[31] & x_a[30] & (!x_b[30]));//depth1
 
  assign XOR[29] = x_a[29] ^ (!x_b[29]);
  assign XOR[28] = x_a[28] ^ (!x_b[28]);
  assign GT2_15 = (x_a[29] & (!x_b[29])) ^ (XOR[29] & x_a[28] & (!x_b[28]));//depth1
  
  assign temp[8] = XOR[31] & XOR[30] & GT2_15;//depth2
  assign GT4_8 = temp[8] ^ GT2_16;//depth2
  ///////////////////////////////////////////// 
  assign XOR[27]= x_a[27] ^ (!x_b[27]);
  assign XOR[26]= x_a[26] ^ (!x_b[26]);
  assign GT2_14 = (x_a[27] & (!x_b[27])) ^ (XOR[27] & x_a[26] & (!x_b[26]));//depth1
 
  assign XOR[25] = x_a[25] ^ (!x_b[25]);
  assign XOR[24] = x_a[24] ^ (!x_b[24]);
  assign GT2_13 = (x_a[25] & (!x_b[25])) ^ (XOR[25] & x_a[24] & (!x_b[24]));//depth1
  
  //assign temp[7] = XOR[27] & XOR[26] & GT2_13;//depth2
  //assign GT4_7 = temp[7] ^ GT2_14;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[12]= XOR[31] & XOR[30] & XOR[29] & XOR[28];//depth1
  assign AND31_28= (temp[12] & GT2_14) ^ (temp[12] & XOR[27] & XOR[26] & GT2_13);//depth2
  assign GT8_4 = AND31_28 ^ GT4_8;
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[23]= x_a[23] ^ (!x_b[23]);
  assign XOR[22]= x_a[22] ^ (!x_b[22]);
  assign GT2_12 = (x_a[23] & (!x_b[23])) ^ (XOR[23] & x_a[22] & (!x_b[22])); //depth1
 
  assign XOR[21] = x_a[21] ^ (!x_b[21]);
  assign XOR[20] = x_a[20] ^ (!x_b[20]);
  assign GT2_11 = (x_a[21] & (!x_b[21])) ^ (XOR[21] & x_a[20] & (!x_b[20])); //depth1
  
  assign temp[6] = XOR[23] & XOR[22] & GT2_11;//depth2
  assign GT4_6 = temp[6] ^ GT2_12;//depth2
  ///////////////////////////////////////////// 
  assign XOR[19]= x_a[19] ^ (!x_b[19]);
  assign XOR[18]= x_a[18] ^ (!x_b[18]);
  assign GT2_10 = (x_a[19] & (!x_b[19])) ^ (XOR[19] & x_a[18] & (!x_b[18]));//depth1
 
  assign XOR[17] = x_a[17] ^ (!x_b[17]);
  assign XOR[16] = x_a[16] ^ (!x_b[16]);
  assign GT2_9 = (x_a[17] & (!x_b[17])) ^ (XOR[17] & x_a[16] & (!x_b[16]));//depth1
  
  //assign temp[5] = XOR[19] & XOR[18] & GT2_9;//depth2
  //assign GT4_5 = temp[5] ^ GT2_10;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[11]= XOR[23] & XOR[22] & XOR[21] & XOR[20];//depth1
  assign AND23_20= (temp[11] & GT2_10) ^ (temp[11] & XOR[19] & XOR[18] & GT2_9);//depth2
  assign GT8_3 = AND23_20 ^ GT4_6;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign AND27_24= XOR[27] & XOR[26] & XOR[25] & XOR[24];//depth1
  assign temp[14]= AND27_24& temp[12];//depth2
  assign AND31_24=temp[14]&GT8_3;//depth3
  assign GT16_2 = AND31_24 ^ GT8_4;//depth3
  /////////////////////////////////////////////
  /////////////////////////////////////////////
  ////////////////////////////////////////////
  assign XOR[15]= x_a[15] ^ (!x_b[15]); //depth1
  assign XOR[14]= x_a[14] ^ (!x_b[14]);
  assign GT2_8 = (x_a[15] & (!x_b[15])) ^ (XOR[15] & x_a[14] & (!x_b[14]));//depth1
 
  assign XOR[13] = x_a[13] ^ (!x_b[13]);
  assign XOR[12] = x_a[12] ^ (!x_b[12]);
  assign GT2_7 = (x_a[13] & (!x_b[13])) ^ (XOR[13] & x_a[12] & (!x_b[12]));//depth1
  
  assign temp[4] = XOR[15] & XOR[14] & GT2_7;//depth2
  assign GT4_4 = temp[4] ^ GT2_8;//depth2
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[11]= x_a[11] ^ (!x_b[11]);
  assign XOR[10]= x_a[10] ^ (!x_b[10]);
  assign GT2_6 = (x_a[11] & (!x_b[11])) ^ (XOR[11] & x_a[10] & (!x_b[10]));//depth1
 
  assign XOR[9] = x_a[9] ^ (!x_b[9]);
  assign XOR[8] = x_a[8] ^ (!x_b[8]);
  assign GT2_5 = (x_a[9] & (!x_b[9])) ^ (XOR[9] & x_a[8] & (!x_b[8]));//depth1
  
  //assign temp[3] = XOR[11] & XOR[10] & GT2_5;//depth2
  //assign GT4_3 = temp[3] ^ GT2_6;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[10]= XOR[15] & XOR[14] & XOR[13] & XOR[12];//depth1
  assign AND15_12= (temp[10] & GT2_6) ^ (temp[10] & XOR[11] & XOR[10] & GT2_5);//depth2
  assign GT8_2 = AND15_12 ^ GT4_4;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[7]= x_a[7] ^ (!x_b[7]);
  assign XOR[6]= x_a[6] ^ (!x_b[6]);
  assign GT2_4 = (x_a[7] & (!x_b[7])) ^ (XOR[7] & x_a[6] & (!x_b[6]));//depth1
 
  assign XOR[5] = x_a[5] ^ (!x_b[5]);
  assign XOR[4] = x_a[4] ^ (!x_b[4]);
  assign GT2_3  = (x_a[5] & (!x_b[5])) ^ (XOR[5] & x_a[4] & (!x_b[4]));//depth1
  
  assign temp[2] = XOR[7] & XOR[6] & GT2_3;//depth2
  assign GT4_2 = temp[2] ^ GT2_4;//depth2
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[3]= x_a[3] ^ (!x_b[3]);
  assign XOR[2]= x_a[2] ^ (!x_b[2]);
  assign GT2_2 = (x_a[3] & (!x_b[3])) ^ (XOR[3] & x_a[2] & (!x_b[2]));//depth1
 
  assign XOR[1] = x_a[1] ^ (!x_b[1]);
  assign XOR[0] = x_a[0] ^ (!x_b[0]);
  assign GT2_1  = (x_a[1] & (!x_b[1])) ^ (XOR[1] & x_a[0] & (!x_b[0]));//depth1
  
  //assign temp[1] = XOR[3] & XOR[2] & GT2_1;//depth2
  //assign GT4_1 = temp[1] ^ GT2_2;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[9]= XOR[7] & XOR[6] & XOR[5] & XOR[4];//depth1
  assign AND7_4= (temp[9] & GT2_2) ^ (temp[9] & XOR[3] & XOR[2] & GT2_1);//depth2
  assign GT8_1 = AND7_4 ^ GT4_2;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign AND11_8= XOR[11] & XOR[10] & XOR[9] & XOR[8];//depth1
  assign temp[13]= AND11_8& temp[10];//depth2
  //assign XOR15_8=temp[13]&GT8_1;//depth3
  //assign GT16_1 = XOR15_8 ^ GT8_2;//depth3
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign AND19_16= XOR[19] & XOR[18] & XOR[17] & XOR[16];//depth1
  assign temp[15]= AND19_16& AND27_24& temp[12]&temp[11];//depth2
  assign AND31_16= (temp[15]&temp[13]&GT8_1) ^ (temp[15]& GT8_2);//depth3
  assign GT32_1 = AND31_16 ^ GT16_2;//depth3
   /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////

  assign wx = GT32_1;
endmodule



