module main(input wire a, output wire b);
   assign b = a;
endmodule // main
