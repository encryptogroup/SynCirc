module main(input wire a, output wire b);
   assign b = 0;
endmodule // main
