module COMP8 (x_a, x_b, wx);
  input  [7:0] x_a, x_b;
  output wx;
  wire [7:0] XOR;
  wire [3:0] temp;
  wire GT2_4,GT2_3,GT2_2,GT2_1;
  wire GT4_2,GT4_1;
  wire GT8_1;
  wire AND7_4; 
  
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[7]= x_a[7] ^ (!x_b[7]);
  assign XOR[6]= x_a[6] ^ (!x_b[6]);
  assign GT2_4 = (x_a[7] & (!x_b[7])) ^ (XOR[7] & x_a[6] & (!x_b[6]));//depth1
 
  assign XOR[5] = x_a[5] ^ (!x_b[5]);
  assign XOR[4] = x_a[4] ^ (!x_b[4]);
  assign GT2_3  = (x_a[5] & (!x_b[5])) ^ (XOR[5] & x_a[4] & (!x_b[4]));//depth1
  
  assign temp[2] = XOR[7] & XOR[6] & GT2_3;//depth2
  assign GT4_2 = temp[2] ^ GT2_4;//depth2
  /////////////////////////////////////////////////////////////////////////////
  assign XOR[3]= x_a[3] ^ (!x_b[3]);
  assign XOR[2]= x_a[2] ^ (!x_b[2]);
  assign GT2_2 = (x_a[3] & (!x_b[3])) ^ (XOR[3] & x_a[2] & (!x_b[2]));//depth1
 
  assign XOR[1] = x_a[1] ^ (!x_b[1]);
  assign XOR[0] = x_a[0] ^ (!x_b[0]);
  assign GT2_1  = (x_a[1] & (!x_b[1])) ^ (XOR[1] & x_a[0] & (!x_b[0]));//depth1
  
  //assign temp[1] = XOR[3] & XOR[2] & GT2_1;//depth2
  //assign GT4_1 = temp[1] ^ GT2_2;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////
  assign temp[3]= XOR[7] & XOR[6] & XOR[5] & XOR[4];//depth1
  assign AND7_4= (temp[3] & GT2_2) ^ (temp[3] & XOR[3] & XOR[2] & GT2_1);//depth2
  assign GT8_1 = AND7_4 ^ GT4_2;//depth2
  /////////////////////////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////////////////////////


  assign wx = GT8_1;
endmodule



